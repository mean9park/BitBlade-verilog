`timescale 1ns / 1ps

// Have to packing data from all the Processing element!!!! 
// So only one wire_packing is used in bitblade_column.v

module Weight_Wire_packing(
    input clk,
    input reset,
    
    input [31:0] sorted_weight_1, sorted_weight_2, sorted_weight_3, sorted_weight_4, sorted_weight_5, sorted_weight_6, sorted_weight_7, sorted_weight_8, 
    sorted_weight_9, sorted_weight_10, sorted_weight_11, sorted_weight_12, sorted_weight_13, sorted_weight_14, sorted_weight_15, sorted_weight_16, 

    output [31:0] packed_weight_1, packed_weight_2, packed_weight_3, packed_weight_4, packed_weight_5, packed_weight_6, packed_weight_7, packed_weight_8, 
    packed_weight_9, packed_weight_10, packed_weight_11, packed_weight_12, packed_weight_13, packed_weight_14, packed_weight_15, packed_weight_16
);
    
    assign packed_weight_1 = {sorted_weight_16[1:0], sorted_weight_15[1:0], sorted_weight_14[1:0], sorted_weight_13[1:0], sorted_weight_12[1:0], sorted_weight_11[1:0], sorted_weight_10[1:0], sorted_weight_9[1:0], sorted_weight_8[1:0], sorted_weight_7[1:0], sorted_weight_6[1:0], sorted_weight_5[1:0], sorted_weight_4[1:0], sorted_weight_3[1:0], sorted_weight_2[1:0], sorted_weight_1[1:0]};
    assign packed_weight_2 = {sorted_weight_16[3:2], sorted_weight_15[3:2], sorted_weight_14[3:2], sorted_weight_13[3:2], sorted_weight_12[3:2], sorted_weight_11[3:2], sorted_weight_10[3:2], sorted_weight_9[3:2], sorted_weight_8[3:2], sorted_weight_7[3:2], sorted_weight_6[3:2], sorted_weight_5[3:2], sorted_weight_4[3:2], sorted_weight_3[3:2], sorted_weight_2[3:2], sorted_weight_1[3:2]};
    assign packed_weight_3 = {sorted_weight_16[5:4], sorted_weight_15[5:4], sorted_weight_14[5:4], sorted_weight_13[5:4], sorted_weight_12[5:4], sorted_weight_11[5:4], sorted_weight_10[5:4], sorted_weight_9[5:4], sorted_weight_8[5:4], sorted_weight_7[5:4], sorted_weight_6[5:4], sorted_weight_5[5:4], sorted_weight_4[5:4], sorted_weight_3[5:4], sorted_weight_2[5:4], sorted_weight_1[5:4]};
    assign packed_weight_4 = {sorted_weight_16[7:6], sorted_weight_15[7:6], sorted_weight_14[7:6], sorted_weight_13[7:6], sorted_weight_12[7:6], sorted_weight_11[7:6], sorted_weight_10[7:6], sorted_weight_9[7:6], sorted_weight_8[7:6], sorted_weight_7[7:6], sorted_weight_6[7:6], sorted_weight_5[7:6], sorted_weight_4[7:6], sorted_weight_3[7:6], sorted_weight_2[7:6], sorted_weight_1[7:6]};
    assign packed_weight_5 = {sorted_weight_16[9:8], sorted_weight_15[9:8], sorted_weight_14[9:8], sorted_weight_13[9:8], sorted_weight_12[9:8], sorted_weight_11[9:8], sorted_weight_10[9:8], sorted_weight_9[9:8], sorted_weight_8[9:8], sorted_weight_7[9:8], sorted_weight_6[9:8], sorted_weight_5[9:8], sorted_weight_4[9:8], sorted_weight_3[9:8], sorted_weight_2[9:8], sorted_weight_1[9:8]};
    assign packed_weight_6 = {sorted_weight_16[11:10], sorted_weight_15[11:10], sorted_weight_14[11:10], sorted_weight_13[11:10], sorted_weight_12[11:10], sorted_weight_11[11:10], sorted_weight_10[11:10], sorted_weight_9[11:10], sorted_weight_8[11:10], sorted_weight_7[11:10], sorted_weight_6[11:10], sorted_weight_5[11:10], sorted_weight_4[11:10], sorted_weight_3[11:10], sorted_weight_2[11:10], sorted_weight_1[11:10]};
    assign packed_weight_7 = {sorted_weight_16[13:12], sorted_weight_15[13:12], sorted_weight_14[13:12], sorted_weight_13[13:12], sorted_weight_12[13:12], sorted_weight_11[13:12], sorted_weight_10[13:12], sorted_weight_9[13:12], sorted_weight_8[13:12], sorted_weight_7[13:12], sorted_weight_6[13:12], sorted_weight_5[13:12], sorted_weight_4[13:12], sorted_weight_3[13:12], sorted_weight_2[13:12], sorted_weight_1[13:12]};
    assign packed_weight_8 = {sorted_weight_16[15:14], sorted_weight_15[15:14], sorted_weight_14[15:14], sorted_weight_13[15:14], sorted_weight_12[15:14], sorted_weight_11[15:14], sorted_weight_10[15:14], sorted_weight_9[15:14], sorted_weight_8[15:14], sorted_weight_7[15:14], sorted_weight_6[15:14], sorted_weight_5[15:14], sorted_weight_4[15:14], sorted_weight_3[15:14], sorted_weight_2[15:14], sorted_weight_1[15:14]};
    assign packed_weight_9 = {sorted_weight_16[17:16], sorted_weight_15[17:16], sorted_weight_14[17:16], sorted_weight_13[17:16], sorted_weight_12[17:16], sorted_weight_11[17:16], sorted_weight_10[17:16], sorted_weight_9[17:16], sorted_weight_8[17:16], sorted_weight_7[17:16], sorted_weight_6[17:16], sorted_weight_5[17:16], sorted_weight_4[17:16], sorted_weight_3[17:16], sorted_weight_2[17:16], sorted_weight_1[17:16]};
    assign packed_weight_10 = {sorted_weight_16[19:18], sorted_weight_15[19:18], sorted_weight_14[19:18], sorted_weight_13[19:18], sorted_weight_12[19:18], sorted_weight_11[19:18], sorted_weight_10[19:18], sorted_weight_9[19:18], sorted_weight_8[19:18], sorted_weight_7[19:18], sorted_weight_6[19:18], sorted_weight_5[19:18], sorted_weight_4[19:18], sorted_weight_3[19:18], sorted_weight_2[19:18], sorted_weight_1[19:18]};
    assign packed_weight_11 = {sorted_weight_16[21:20], sorted_weight_15[21:20], sorted_weight_14[21:20], sorted_weight_13[21:20], sorted_weight_12[21:20], sorted_weight_11[21:20], sorted_weight_10[21:20], sorted_weight_9[21:20], sorted_weight_8[21:20], sorted_weight_7[21:20], sorted_weight_6[21:20], sorted_weight_5[21:20], sorted_weight_4[21:20], sorted_weight_3[21:20], sorted_weight_2[21:20], sorted_weight_1[21:20]};
    assign packed_weight_12 = {sorted_weight_16[23:22], sorted_weight_15[23:22], sorted_weight_14[23:22], sorted_weight_13[23:22], sorted_weight_12[23:22], sorted_weight_11[23:22], sorted_weight_10[23:22], sorted_weight_9[23:22], sorted_weight_8[23:22], sorted_weight_7[23:22], sorted_weight_6[23:22], sorted_weight_5[23:22], sorted_weight_4[23:22], sorted_weight_3[23:22], sorted_weight_2[23:22], sorted_weight_1[23:22]};
    assign packed_weight_13 = {sorted_weight_16[25:24], sorted_weight_15[25:24], sorted_weight_14[25:24], sorted_weight_13[25:24], sorted_weight_12[25:24], sorted_weight_11[25:24], sorted_weight_10[25:24], sorted_weight_9[25:24], sorted_weight_8[25:24], sorted_weight_7[25:24], sorted_weight_6[25:24], sorted_weight_5[25:24], sorted_weight_4[25:24], sorted_weight_3[25:24], sorted_weight_2[25:24], sorted_weight_1[25:24]};
    assign packed_weight_14 = {sorted_weight_16[27:26], sorted_weight_15[27:26], sorted_weight_14[27:26], sorted_weight_13[27:26], sorted_weight_12[27:26], sorted_weight_11[27:26], sorted_weight_10[27:26], sorted_weight_9[27:26], sorted_weight_8[27:26], sorted_weight_7[27:26], sorted_weight_6[27:26], sorted_weight_5[27:26], sorted_weight_4[27:26], sorted_weight_3[27:26], sorted_weight_2[27:26], sorted_weight_1[27:26]};
    assign packed_weight_15 = {sorted_weight_16[29:28], sorted_weight_15[29:28], sorted_weight_14[29:28], sorted_weight_13[29:28], sorted_weight_12[29:28], sorted_weight_11[29:28], sorted_weight_10[29:28], sorted_weight_9[29:28], sorted_weight_8[29:28], sorted_weight_7[29:28], sorted_weight_6[29:28], sorted_weight_5[29:28], sorted_weight_4[29:28], sorted_weight_3[29:28], sorted_weight_2[29:28], sorted_weight_1[29:28]};
    assign packed_weight_16 = {sorted_weight_16[31:30], sorted_weight_15[31:30], sorted_weight_14[31:30], sorted_weight_13[31:30], sorted_weight_12[31:30], sorted_weight_11[31:30], sorted_weight_10[31:30], sorted_weight_9[31:30], sorted_weight_8[31:30], sorted_weight_7[31:30], sorted_weight_6[31:30], sorted_weight_5[31:30], sorted_weight_4[31:30], sorted_weight_3[31:30], sorted_weight_2[31:30], sorted_weight_1[31:30]};

endmodule