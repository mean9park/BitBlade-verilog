`timescale 1ns / 1ps

// I have two seperate file for input, weight 
// But they are the same!

module Input_Wire_packing(
    input clk,
    input reset,
    
    input [31:0] sorted_input_1, sorted_input_2, sorted_input_3, sorted_input_4, sorted_input_5, sorted_input_6, sorted_input_7, sorted_input_8, 
    sorted_input_9, sorted_input_10, sorted_input_11, sorted_input_12, sorted_input_13, sorted_input_14, sorted_input_15, sorted_input_16, 

    output [31:0] packed_input_1, packed_input_2, packed_input_3, packed_input_4, packed_input_5, packed_input_6, packed_input_7, packed_input_8, 
    packed_input_9, packed_input_10, packed_input_11, packed_input_12, packed_input_13, packed_input_14, packed_input_15, packed_input_16
);
    
    assign packed_input_1 = {sorted_input_16[1:0], sorted_input_15[1:0], sorted_input_14[1:0], sorted_input_13[1:0], sorted_input_12[1:0], sorted_input_11[1:0], sorted_input_10[1:0], sorted_input_9[1:0], sorted_input_8[1:0], sorted_input_7[1:0], sorted_input_6[1:0], sorted_input_5[1:0], sorted_input_4[1:0], sorted_input_3[1:0], sorted_input_2[1:0], sorted_input_1[1:0]};
    assign packed_input_2 = {sorted_input_16[3:2], sorted_input_15[3:2], sorted_input_14[3:2], sorted_input_13[3:2], sorted_input_12[3:2], sorted_input_11[3:2], sorted_input_10[3:2], sorted_input_9[3:2], sorted_input_8[3:2], sorted_input_7[3:2], sorted_input_6[3:2], sorted_input_5[3:2], sorted_input_4[3:2], sorted_input_3[3:2], sorted_input_2[3:2], sorted_input_1[3:2]};
    assign packed_input_3 = {sorted_input_16[5:4], sorted_input_15[5:4], sorted_input_14[5:4], sorted_input_13[5:4], sorted_input_12[5:4], sorted_input_11[5:4], sorted_input_10[5:4], sorted_input_9[5:4], sorted_input_8[5:4], sorted_input_7[5:4], sorted_input_6[5:4], sorted_input_5[5:4], sorted_input_4[5:4], sorted_input_3[5:4], sorted_input_2[5:4], sorted_input_1[5:4]};
    assign packed_input_4 = {sorted_input_16[7:6], sorted_input_15[7:6], sorted_input_14[7:6], sorted_input_13[7:6], sorted_input_12[7:6], sorted_input_11[7:6], sorted_input_10[7:6], sorted_input_9[7:6], sorted_input_8[7:6], sorted_input_7[7:6], sorted_input_6[7:6], sorted_input_5[7:6], sorted_input_4[7:6], sorted_input_3[7:6], sorted_input_2[7:6], sorted_input_1[7:6]};
    assign packed_input_5 = {sorted_input_16[9:8], sorted_input_15[9:8], sorted_input_14[9:8], sorted_input_13[9:8], sorted_input_12[9:8], sorted_input_11[9:8], sorted_input_10[9:8], sorted_input_9[9:8], sorted_input_8[9:8], sorted_input_7[9:8], sorted_input_6[9:8], sorted_input_5[9:8], sorted_input_4[9:8], sorted_input_3[9:8], sorted_input_2[9:8], sorted_input_1[9:8]};
    assign packed_input_6 = {sorted_input_16[11:10], sorted_input_15[11:10], sorted_input_14[11:10], sorted_input_13[11:10], sorted_input_12[11:10], sorted_input_11[11:10], sorted_input_10[11:10], sorted_input_9[11:10], sorted_input_8[11:10], sorted_input_7[11:10], sorted_input_6[11:10], sorted_input_5[11:10], sorted_input_4[11:10], sorted_input_3[11:10], sorted_input_2[11:10], sorted_input_1[11:10]};
    assign packed_input_7 = {sorted_input_16[13:12], sorted_input_15[13:12], sorted_input_14[13:12], sorted_input_13[13:12], sorted_input_12[13:12], sorted_input_11[13:12], sorted_input_10[13:12], sorted_input_9[13:12], sorted_input_8[13:12], sorted_input_7[13:12], sorted_input_6[13:12], sorted_input_5[13:12], sorted_input_4[13:12], sorted_input_3[13:12], sorted_input_2[13:12], sorted_input_1[13:12]};
    assign packed_input_8 = {sorted_input_16[15:14], sorted_input_15[15:14], sorted_input_14[15:14], sorted_input_13[15:14], sorted_input_12[15:14], sorted_input_11[15:14], sorted_input_10[15:14], sorted_input_9[15:14], sorted_input_8[15:14], sorted_input_7[15:14], sorted_input_6[15:14], sorted_input_5[15:14], sorted_input_4[15:14], sorted_input_3[15:14], sorted_input_2[15:14], sorted_input_1[15:14]};
    assign packed_input_9 = {sorted_input_16[17:16], sorted_input_15[17:16], sorted_input_14[17:16], sorted_input_13[17:16], sorted_input_12[17:16], sorted_input_11[17:16], sorted_input_10[17:16], sorted_input_9[17:16], sorted_input_8[17:16], sorted_input_7[17:16], sorted_input_6[17:16], sorted_input_5[17:16], sorted_input_4[17:16], sorted_input_3[17:16], sorted_input_2[17:16], sorted_input_1[17:16]};
    assign packed_input_10 = {sorted_input_16[19:18], sorted_input_15[19:18], sorted_input_14[19:18], sorted_input_13[19:18], sorted_input_12[19:18], sorted_input_11[19:18], sorted_input_10[19:18], sorted_input_9[19:18], sorted_input_8[19:18], sorted_input_7[19:18], sorted_input_6[19:18], sorted_input_5[19:18], sorted_input_4[19:18], sorted_input_3[19:18], sorted_input_2[19:18], sorted_input_1[19:18]};
    assign packed_input_11 = {sorted_input_16[21:20], sorted_input_15[21:20], sorted_input_14[21:20], sorted_input_13[21:20], sorted_input_12[21:20], sorted_input_11[21:20], sorted_input_10[21:20], sorted_input_9[21:20], sorted_input_8[21:20], sorted_input_7[21:20], sorted_input_6[21:20], sorted_input_5[21:20], sorted_input_4[21:20], sorted_input_3[21:20], sorted_input_2[21:20], sorted_input_1[21:20]};
    assign packed_input_12 = {sorted_input_16[23:22], sorted_input_15[23:22], sorted_input_14[23:22], sorted_input_13[23:22], sorted_input_12[23:22], sorted_input_11[23:22], sorted_input_10[23:22], sorted_input_9[23:22], sorted_input_8[23:22], sorted_input_7[23:22], sorted_input_6[23:22], sorted_input_5[23:22], sorted_input_4[23:22], sorted_input_3[23:22], sorted_input_2[23:22], sorted_input_1[23:22]};
    assign packed_input_13 = {sorted_input_16[25:24], sorted_input_15[25:24], sorted_input_14[25:24], sorted_input_13[25:24], sorted_input_12[25:24], sorted_input_11[25:24], sorted_input_10[25:24], sorted_input_9[25:24], sorted_input_8[25:24], sorted_input_7[25:24], sorted_input_6[25:24], sorted_input_5[25:24], sorted_input_4[25:24], sorted_input_3[25:24], sorted_input_2[25:24], sorted_input_1[25:24]};
    assign packed_input_14 = {sorted_input_16[27:26], sorted_input_15[27:26], sorted_input_14[27:26], sorted_input_13[27:26], sorted_input_12[27:26], sorted_input_11[27:26], sorted_input_10[27:26], sorted_input_9[27:26], sorted_input_8[27:26], sorted_input_7[27:26], sorted_input_6[27:26], sorted_input_5[27:26], sorted_input_4[27:26], sorted_input_3[27:26], sorted_input_2[27:26], sorted_input_1[27:26]};
    assign packed_input_15 = {sorted_input_16[29:28], sorted_input_15[29:28], sorted_input_14[29:28], sorted_input_13[29:28], sorted_input_12[29:28], sorted_input_11[29:28], sorted_input_10[29:28], sorted_input_9[29:28], sorted_input_8[29:28], sorted_input_7[29:28], sorted_input_6[29:28], sorted_input_5[29:28], sorted_input_4[29:28], sorted_input_3[29:28], sorted_input_2[29:28], sorted_input_1[29:28]};
    assign packed_input_16 = {sorted_input_16[31:30], sorted_input_15[31:30], sorted_input_14[31:30], sorted_input_13[31:30], sorted_input_12[31:30], sorted_input_11[31:30], sorted_input_10[31:30], sorted_input_9[31:30], sorted_input_8[31:30], sorted_input_7[31:30], sorted_input_6[31:30], sorted_input_5[31:30], sorted_input_4[31:30], sorted_input_3[31:30], sorted_input_2[31:30], sorted_input_1[31:30]};

endmodule